library verilog;
use verilog.vl_types.all;
entity gate_vlg_vec_tst is
end gate_vlg_vec_tst;
