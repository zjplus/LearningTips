library verilog;
use verilog.vl_types.all;
entity FrequencyDivision097_vlg_vec_tst is
end FrequencyDivision097_vlg_vec_tst;
