LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY voter097 IS
PORT(A0,A1,A2,A3,A4:IN STD_LOGIC;
Y:OUT STD_LOGIC);
END ENTITY voter097;

ARCHITECTURE TOUPIAOQI OF voter097 IS
BEGIN PROCESS(A0,A1,A2,A3,A4)
VARIABLE SUM:INTEGER;
BEGIN
SUM:=0;
IF A0='1' THEN SUM:=SUM+1;END IF;
IF A1='1' THEN SUM:=SUM+1;END IF;
IF A2='1' THEN SUM:=SUM+1;END IF;
IF A3='1' THEN SUM:=SUM+1;END IF;
IF A4='1' THEN SUM:=SUM+1;END IF;
IF SUM>2 THEN Y<='1';
ELSE Y<='0';
END IF;
END PROCESS;
END TOUPIAOQI;