library verilog;
use verilog.vl_types.all;
entity FrequencyDivision097 is
    port(
        clk             : in     vl_logic;
        Q1              : inout  vl_logic;
        Q2              : out    vl_logic
    );
end FrequencyDivision097;
