library verilog;
use verilog.vl_types.all;
entity gate097_vlg_vec_tst is
end gate097_vlg_vec_tst;
