library verilog;
use verilog.vl_types.all;
entity gate_vlg_check_tst is
    port(
        e               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end gate_vlg_check_tst;
