library verilog;
use verilog.vl_types.all;
entity FrequencyDivision097_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        Q1              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end FrequencyDivision097_vlg_sample_tst;
