library verilog;
use verilog.vl_types.all;
entity Clock_097_vlg_vec_tst is
end Clock_097_vlg_vec_tst;
