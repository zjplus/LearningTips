library verilog;
use verilog.vl_types.all;
entity counter097_vlg_vec_tst is
end counter097_vlg_vec_tst;
