library verilog;
use verilog.vl_types.all;
entity voter097_vlg_vec_tst is
end voter097_vlg_vec_tst;
