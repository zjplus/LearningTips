library verilog;
use verilog.vl_types.all;
entity Clock_097_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Clock_097_vlg_sample_tst;
